.title KiCad schematic
.include "C:/AE/MAX4719/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/MAX4719/_models/MAX4719.FAM"
R1 /COM1 0 {RCOM1}
V6 /CTRL2 0 PULSE( 0 5 4m 10n 10n 6m 12m ) 
R2 /COM2 0 {RCOM2}
V7 /NC1 0 DC 3 SIN( 3 1 1k 0 0 0 ) AC 1  
V1 VDD 0 DC {VSUPPLY} 
XU1 VDD 0 C2012X7R2A104K125AA_p
XU2 VDD /NO1 /COM1 /CTRL1 /NC1 0 /NC2 /CTRL2 /COM2 /NO2 MAX4719
V2 /NO2 0 DC 2 SIN( 2 1 2k 0 0 0 ) AC 1  
V4 /NO1 0 DC 3 SIN( 3 0.5 2k 0 0 0 ) AC 1  
V3 /CTRL1 0 PULSE( 0 5 6m 10n 10n 4m 8m ) 
V5 /NC2 0 DC 2 SIN( 2 0.5 1k 0 0 0 ) AC 1  
.end
